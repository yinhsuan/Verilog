//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
//0511049

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
wire     [32-1:0] data_o;
assign data_o[15:0] = data_i[15:0] ;
assign data_o[31:16] = data_i[15] ? 16'b1111_1111_1111_1111 : 16'b0000_0000_0000_0000;

//Sign extended
          
endmodule      
     